pBAV       �c      @       �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@             @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               D^
BX�hh^�&^�	��~�N���L��	&�	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                