pBAV       �       @       �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@             @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               V�d N � T6Td l 2� N�Z                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               