pBAV       @�       @       �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@             @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               V�d N � T6Td * 2� N�Z                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               