pBAV       ��     
 @       �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@             @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               N~	`n J��L	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          